`include "Half_Add.sv"  
`include "FetchInstruction.sv"
`include "Registers.sv"
`include "Full_Add.sv"
`include "Controls.sv"
`include "ALU_Control.sv"


  
  






  

	
    